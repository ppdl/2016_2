library verilog;
use verilog.vl_types.all;
entity testbench0 is
end testbench0;
